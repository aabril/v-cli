module main

import commands

fn main() {
    commands.set()
}

